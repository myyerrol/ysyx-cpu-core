module fsm_top(

);



endmodule
