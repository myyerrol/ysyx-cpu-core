`include "Config.v"

module AXI4LiteM(
    input  wire                       iClock,
    input  wire                       iReset,
    input  wire [`MODE_WIDTH - 1 : 0] iMode,
    input  wire [`ADDR_WIDTH - 1 : 0] iAddr,
    input  wire [`DATA_WIDTH - 1 : 0] iData,
    input  wire [`MASK_WIDTH - 1 : 0] iMask,
    input  wire                       iValid,
    output wire [`DATA_WIDTH - 1 : 0] oData,
    output wire [`RESP_WIDTH - 1 : 0] oResp,

    input  wire                       pAXI4_ar_ready,
    output wire                       pAXI4_ar_valid,
    output wire [`ADDR_WIDTH - 1 : 0] pAXI4_ar_bits_addr,

    input  wire                       pAXI4_r_valid,
    input  wire [`DATA_WIDTH - 1 : 0] pAXI4_r_bits_data,
    input  wire [`RESP_WIDTH - 1 : 0] pAXI4_r_bits_resp,
    output wire                       pAXI4_r_ready,

    input  wire                       pAXI4_aw_ready,
    output wire                       pAXI4_aw_valid,
    output wire [`ADDR_WIDTH - 1 : 0] pAXI4_aw_bits_addr,

    input  wire                       pAXI4_w_ready,
    output wire                       pAXI4_w_valid,
    output wire [`DATA_WIDTH - 1 : 0] pAXI4_w_bits_data,
    output wire [`MASK_WIDTH - 1 : 0] pAXI4_w_bits_strb,

    input  wire                       pAXI4_b_valid,
    input  wire [`RESP_WIDTH - 1 : 0] pAXI4_b_bits_resp,
    output wire                       pAXI4_b_ready
);

    always @(posedge iClock) begin
`ifdef VTRACE_MONITOR
        $display("[vtrace] clock:      %d, reset:      %d", iClock, iReset);
        $display("[vtrace] state curr: %d, state next: %d", r_state_rd_curr,
                                                            r_state_rd_next);
        $display("[vtrace] arvalid:    %d, arready:    %d, araddr: %x",
                 pAXI4_ar_valid,
                 pAXI4_ar_ready,
                 pAXI4_ar_bits_addr);
        $display("[vtrace] rvalid:     %d, rready:     %d, rdata:  %x, rresp: %d",
                 pAXI4_r_valid,
                 pAXI4_r_ready,
                 oData,
                 pAXI4_r_bits_resp);
`endif
    end

    //-------------------------------------------------------------------------
    parameter P_STATE_IDLE     = 'd0;
    parameter P_STATE_RD_TRANS = 'd1;
    parameter P_STATE_RD_END   = 'd2;

    reg [2 : 0] r_state_rd_curr;
    reg [2 : 0] r_state_rd_next;

    //-------------------------------------------------------------------------
    wire                       w_arvalid;
    wire [`ADDR_WIDTH - 1 : 0] w_araddr;
    wire [`DATA_WIDTH - 1 : 0] w_ardata;

    wire                       w_rd_start;
    wire                       w_rd_last;
    wire                       w_rd_addr_handshake;
    wire                       w_rd_data_handshake;

    //-------------------------------------------------------------------------
    reg                       r_rready;
    reg [`ADDR_WIDTH - 1 : 0] r_araddr;
    reg [`DATA_WIDTH - 1 : 0] r_rdata;

    reg                       r_awvalid;
    reg [`ADDR_WIDTH - 1 : 0] r_awaddr;
    reg                       r_wvalid;
    reg [`DATA_WIDTH - 1 : 0] r_wdata;
    reg [`MASK_WIDTH - 1 : 0] r_wstrb;
    reg                       r_bready;

    //-------------------------------------------------------------------------
    assign oData               = (iReset) ? `DATA_WIDTH'b0 : r_rdata;
    assign oResp               = pAXI4_r_bits_resp;

    assign pAXI4_ar_valid      = w_arvalid;
    assign pAXI4_ar_bits_addr  = r_araddr;
    assign pAXI4_r_ready       = r_rready;
    assign pAXI4_aw_valid      = r_awvalid;
    assign pAXI4_aw_bits_addr  = r_awaddr;
    assign pAXI4_w_valid       = r_wvalid;
    assign pAXI4_w_bits_data   = r_wdata;
    assign pAXI4_w_bits_strb   = r_wstrb;
    assign pAXI4_b_ready       = 1'b1;

    assign w_arvalid           = iValid;
    assign w_araddr            = (iReset) ? `ADDR_WIDTH'b0 : iAddr;

    assign w_rd_start          = iValid;
    assign w_rd_last           = r_rready;
    assign w_rd_addr_handshake = pAXI4_ar_valid && pAXI4_ar_ready;
    assign w_rd_data_handshake = pAXI4_r_valid  && pAXI4_r_ready;

    //-------------------------------------------------------------------------
    always @(posedge iClock) begin
        if (iReset) begin
            r_araddr <= `ADDR_WIDTH'b0;
        end
        else if (w_rd_addr_handshake) begin
            r_araddr <= iAddr;
        end
        else begin
            r_araddr <= r_araddr;
        end
    end

    always @(posedge iClock) begin
        if (iReset) begin
            r_rready <= 1'b0;
        end
        else if (w_rd_addr_handshake) begin
            r_rready <= 1'b1;
        end
        else if (w_rd_last) begin
            r_rready <= 1'b0;
        end
        else begin
            r_rready <= r_rready;
        end
    end

    always @(posedge iClock) begin
        if (iReset) begin
            r_rdata <= `DATA_WIDTH'b0;
        end
        else if (w_rd_data_handshake) begin
            r_rdata <= pAXI4_r_bits_data;
        end
        else begin
            r_rdata <= r_rdata;
        end
    end

    //-------------------------------------------------------------------------
    always @(posedge iClock) begin
        if (iReset) begin
            r_state_rd_curr <= P_STATE_IDLE;
        end
        else begin
            r_state_rd_curr <= r_state_rd_next;
        end
    end

    always @(*) begin
        case (r_state_rd_curr)
            P_STATE_IDLE: begin
                if (w_rd_start) begin
                    r_state_rd_next = P_STATE_RD_TRANS;
                end
                else begin
                    r_state_rd_next = P_STATE_IDLE;
                end
            end
            P_STATE_RD_TRANS: begin
                if (w_rd_last) begin
                    r_state_rd_next = P_STATE_RD_END;
                end
                else begin
                    r_state_rd_next = P_STATE_RD_TRANS;
                end
            end
            P_STATE_RD_END: begin
                r_state_rd_next = P_STATE_IDLE;
            end
            default: begin
                r_state_rd_next = P_STATE_IDLE;
            end
        endcase
    end
endmodule
